
module ControlUnity (input clk, reset);



endmodule